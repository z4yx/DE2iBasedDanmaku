// de2i_150_qsys.v

// Generated using ACDS version 15.1 185

`timescale 1 ps / 1 ps
module de2i_150_qsys (
		output wire        altpll_sdram_clk,                              //                     altpll_sdram.clk
		input  wire [3:0]  button_external_connection_export,             //       button_external_connection.export
		output wire        chip_sel_export,                               //                         chip_sel.export
		input  wire        clk_clk,                                       //                              clk.clk
		output wire [0:0]  flash_ssram_tri_state_bridge_out_ssram1_cs_n,  // flash_ssram_tri_state_bridge_out.ssram1_cs_n
		output wire [0:0]  flash_ssram_tri_state_bridge_out_ssram_adsc_n, //                                 .ssram_adsc_n
		output wire [0:0]  flash_ssram_tri_state_bridge_out_ssram_we_n,   //                                 .ssram_we_n
		output wire [0:0]  flash_ssram_tri_state_bridge_out_ssram_oe_n,   //                                 .ssram_oe_n
		inout  wire [31:0] flash_ssram_tri_state_bridge_out_fs_data,      //                                 .fs_data
		output wire [3:0]  flash_ssram_tri_state_bridge_out_ssram_be_n,   //                                 .ssram_be_n
		output wire [0:0]  flash_ssram_tri_state_bridge_out_ssram0_cs_n,  //                                 .ssram0_cs_n
		output wire [21:0] flash_ssram_tri_state_bridge_out_fs_addr,      //                                 .fs_addr
		input  wire [31:0] height_external_connection_export,             //       height_external_connection.export
		output wire [3:0]  led_external_connection_export,                //          led_external_connection.export
		input  wire        mem_master_control_fixed_location,             //               mem_master_control.fixed_location
		input  wire [31:0] mem_master_control_read_base,                  //                                 .read_base
		input  wire [31:0] mem_master_control_read_length,                //                                 .read_length
		input  wire        mem_master_control_go,                         //                                 .go
		output wire        mem_master_control_done,                       //                                 .done
		output wire        mem_master_control_early_done,                 //                                 .early_done
		input  wire        mem_master_user_read_buffer,                   //                  mem_master_user.read_buffer
		output wire [31:0] mem_master_user_buffer_output_data,            //                                 .buffer_output_data
		output wire        mem_master_user_data_available,                //                                 .data_available
		output wire        pcie_clk_clk,                                  //                         pcie_clk.clk
		output wire        pcie_ip_clocks_sim_clk250_export,              //               pcie_ip_clocks_sim.clk250_export
		output wire        pcie_ip_clocks_sim_clk500_export,              //                                 .clk500_export
		output wire        pcie_ip_clocks_sim_clk125_export,              //                                 .clk125_export
		input  wire        pcie_ip_pcie_rstn_export,                      //                pcie_ip_pcie_rstn.export
		input  wire        pcie_ip_pipe_ext_pipe_mode,                    //                 pcie_ip_pipe_ext.pipe_mode
		input  wire        pcie_ip_pipe_ext_phystatus_ext,                //                                 .phystatus_ext
		output wire        pcie_ip_pipe_ext_rate_ext,                     //                                 .rate_ext
		output wire [1:0]  pcie_ip_pipe_ext_powerdown_ext,                //                                 .powerdown_ext
		output wire        pcie_ip_pipe_ext_txdetectrx_ext,               //                                 .txdetectrx_ext
		input  wire        pcie_ip_pipe_ext_rxelecidle0_ext,              //                                 .rxelecidle0_ext
		input  wire [7:0]  pcie_ip_pipe_ext_rxdata0_ext,                  //                                 .rxdata0_ext
		input  wire [2:0]  pcie_ip_pipe_ext_rxstatus0_ext,                //                                 .rxstatus0_ext
		input  wire        pcie_ip_pipe_ext_rxvalid0_ext,                 //                                 .rxvalid0_ext
		input  wire        pcie_ip_pipe_ext_rxdatak0_ext,                 //                                 .rxdatak0_ext
		output wire [7:0]  pcie_ip_pipe_ext_txdata0_ext,                  //                                 .txdata0_ext
		output wire        pcie_ip_pipe_ext_txdatak0_ext,                 //                                 .txdatak0_ext
		output wire        pcie_ip_pipe_ext_rxpolarity0_ext,              //                                 .rxpolarity0_ext
		output wire        pcie_ip_pipe_ext_txcompl0_ext,                 //                                 .txcompl0_ext
		output wire        pcie_ip_pipe_ext_txelecidle0_ext,              //                                 .txelecidle0_ext
		input  wire        pcie_ip_reconfig_busy_busy_altgxb_reconfig,    //            pcie_ip_reconfig_busy.busy_altgxb_reconfig
		output wire [4:0]  pcie_ip_reconfig_fromgxb_0_data,               //       pcie_ip_reconfig_fromgxb_0.data
		input  wire [3:0]  pcie_ip_reconfig_togxb_data,                   //           pcie_ip_reconfig_togxb.data
		input  wire        pcie_ip_refclk_export,                         //                   pcie_ip_refclk.export
		input  wire        pcie_ip_rx_in_rx_datain_0,                     //                    pcie_ip_rx_in.rx_datain_0
		input  wire [39:0] pcie_ip_test_in_test_in,                       //                  pcie_ip_test_in.test_in
		output wire        pcie_ip_tx_out_tx_dataout_0,                   //                   pcie_ip_tx_out.tx_dataout_0
		output wire        pcie_rst_n_reset_n,                            //                       pcie_rst_n.reset_n
		output wire [31:0] pio_size_external_connection_export,           //     pio_size_external_connection.export
		input  wire        reset_reset_n,                                 //                            reset.reset_n
		output wire [12:0] sdram_addr,                                    //                            sdram.addr
		output wire [1:0]  sdram_ba,                                      //                                 .ba
		output wire        sdram_cas_n,                                   //                                 .cas_n
		output wire        sdram_cke,                                     //                                 .cke
		output wire        sdram_cs_n,                                    //                                 .cs_n
		inout  wire [31:0] sdram_dq,                                      //                                 .dq
		output wire [3:0]  sdram_dqm,                                     //                                 .dqm
		output wire        sdram_ras_n,                                   //                                 .ras_n
		output wire        sdram_we_n,                                    //                                 .we_n
		input  wire [31:0] width_external_connection_export               //        width_external_connection.export
	);

	wire         altpll_0_c1_clk;                                    // altpll_0:c1 -> [mm_interconnect_0:altpll_0_c1_clk, rst_controller_002:clk, sram0:clk]
	wire         tristate_conduit_pin_sharer_0_tcm_request;          // tristate_conduit_pin_sharer_0:request -> tristate_conduit_bridge_0:request
	wire  [31:0] tristate_conduit_pin_sharer_0_tcm_fs_data_out;      // tristate_conduit_pin_sharer_0:fs_data -> tristate_conduit_bridge_0:tcs_fs_data
	wire         tristate_conduit_pin_sharer_0_tcm_fs_data_outen;    // tristate_conduit_pin_sharer_0:fs_data_outen -> tristate_conduit_bridge_0:tcs_fs_data_outen
	wire   [0:0] tristate_conduit_pin_sharer_0_tcm_ssram0_cs_n_out;  // tristate_conduit_pin_sharer_0:ssram0_cs_n -> tristate_conduit_bridge_0:tcs_ssram0_cs_n
	wire  [21:0] tristate_conduit_pin_sharer_0_tcm_fs_addr_out;      // tristate_conduit_pin_sharer_0:fs_addr -> tristate_conduit_bridge_0:tcs_fs_addr
	wire   [3:0] tristate_conduit_pin_sharer_0_tcm_ssram_be_n_out;   // tristate_conduit_pin_sharer_0:ssram_be_n -> tristate_conduit_bridge_0:tcs_ssram_be_n
	wire   [0:0] tristate_conduit_pin_sharer_0_tcm_ssram_adsc_n_out; // tristate_conduit_pin_sharer_0:ssram_adsc_n -> tristate_conduit_bridge_0:tcs_ssram_adsc_n
	wire         tristate_conduit_pin_sharer_0_tcm_grant;            // tristate_conduit_bridge_0:grant -> tristate_conduit_pin_sharer_0:grant
	wire   [0:0] tristate_conduit_pin_sharer_0_tcm_ssram1_cs_n_out;  // tristate_conduit_pin_sharer_0:ssram1_cs_n -> tristate_conduit_bridge_0:tcs_ssram1_cs_n
	wire   [0:0] tristate_conduit_pin_sharer_0_tcm_ssram_we_n_out;   // tristate_conduit_pin_sharer_0:ssram_we_n -> tristate_conduit_bridge_0:tcs_ssram_we_n
	wire  [31:0] tristate_conduit_pin_sharer_0_tcm_fs_data_in;       // tristate_conduit_bridge_0:tcs_fs_data_in -> tristate_conduit_pin_sharer_0:fs_data_in
	wire   [0:0] tristate_conduit_pin_sharer_0_tcm_ssram_oe_n_out;   // tristate_conduit_pin_sharer_0:ssram_oe_n -> tristate_conduit_bridge_0:tcs_ssram_oe_n
	wire         ssram0_tcm_data_outen;                              // ssram0:tcm_data_outen -> tristate_conduit_pin_sharer_0:tcs0_data_outen
	wire         ssram0_tcm_outputenable_n_out;                      // ssram0:tcm_outputenable_n_out -> tristate_conduit_pin_sharer_0:tcs0_outputenable_n_out
	wire         ssram0_tcm_request;                                 // ssram0:tcm_request -> tristate_conduit_pin_sharer_0:tcs0_request
	wire   [3:0] ssram0_tcm_byteenable_n_out;                        // ssram0:tcm_byteenable_n_out -> tristate_conduit_pin_sharer_0:tcs0_byteenable_n_out
	wire         ssram0_tcm_write_n_out;                             // ssram0:tcm_write_n_out -> tristate_conduit_pin_sharer_0:tcs0_write_n_out
	wire         ssram0_tcm_begintransfer_n_out;                     // ssram0:tcm_begintransfer_n_out -> tristate_conduit_pin_sharer_0:tcs0_begintransfer_n_out
	wire         ssram0_tcm_grant;                                   // tristate_conduit_pin_sharer_0:tcs0_grant -> ssram0:tcm_grant
	wire         ssram0_tcm_chipselect_n_out;                        // ssram0:tcm_chipselect_n_out -> tristate_conduit_pin_sharer_0:tcs0_chipselect_n_out
	wire  [21:0] ssram0_tcm_address_out;                             // ssram0:tcm_address_out -> tristate_conduit_pin_sharer_0:tcs0_address_out
	wire  [31:0] ssram0_tcm_data_out;                                // ssram0:tcm_data_out -> tristate_conduit_pin_sharer_0:tcs0_data_out
	wire  [31:0] ssram0_tcm_data_in;                                 // tristate_conduit_pin_sharer_0:tcs0_data_in -> ssram0:tcm_data_in
	wire         ssram1_tcm_data_outen;                              // ssram1:tcm_data_outen -> tristate_conduit_pin_sharer_0:tcs1_data_outen
	wire         ssram1_tcm_outputenable_n_out;                      // ssram1:tcm_outputenable_n_out -> tristate_conduit_pin_sharer_0:tcs1_outputenable_n_out
	wire         ssram1_tcm_request;                                 // ssram1:tcm_request -> tristate_conduit_pin_sharer_0:tcs1_request
	wire   [3:0] ssram1_tcm_byteenable_n_out;                        // ssram1:tcm_byteenable_n_out -> tristate_conduit_pin_sharer_0:tcs1_byteenable_n_out
	wire         ssram1_tcm_write_n_out;                             // ssram1:tcm_write_n_out -> tristate_conduit_pin_sharer_0:tcs1_write_n_out
	wire         ssram1_tcm_begintransfer_n_out;                     // ssram1:tcm_begintransfer_n_out -> tristate_conduit_pin_sharer_0:tcs1_begintransfer_n_out
	wire         ssram1_tcm_grant;                                   // tristate_conduit_pin_sharer_0:tcs1_grant -> ssram1:tcm_grant
	wire         ssram1_tcm_chipselect_n_out;                        // ssram1:tcm_chipselect_n_out -> tristate_conduit_pin_sharer_0:tcs1_chipselect_n_out
	wire  [21:0] ssram1_tcm_address_out;                             // ssram1:tcm_address_out -> tristate_conduit_pin_sharer_0:tcs1_address_out
	wire  [31:0] ssram1_tcm_data_out;                                // ssram1:tcm_data_out -> tristate_conduit_pin_sharer_0:tcs1_data_out
	wire  [31:0] ssram1_tcm_data_in;                                 // tristate_conduit_pin_sharer_0:tcs1_data_in -> ssram1:tcm_data_in
	wire  [31:0] mem_master_avalon_master_readdata;                  // mm_interconnect_0:mem_master_avalon_master_readdata -> mem_master:master_readdata
	wire         mem_master_avalon_master_waitrequest;               // mm_interconnect_0:mem_master_avalon_master_waitrequest -> mem_master:master_waitrequest
	wire  [31:0] mem_master_avalon_master_address;                   // mem_master:master_address -> mm_interconnect_0:mem_master_avalon_master_address
	wire         mem_master_avalon_master_read;                      // mem_master:master_read -> mm_interconnect_0:mem_master_avalon_master_read
	wire   [3:0] mem_master_avalon_master_byteenable;                // mem_master:master_byteenable -> mm_interconnect_0:mem_master_avalon_master_byteenable
	wire         mem_master_avalon_master_readdatavalid;             // mm_interconnect_0:mem_master_avalon_master_readdatavalid -> mem_master:master_readdatavalid
	wire   [7:0] mem_master_avalon_master_burstcount;                // mem_master:master_burstcount -> mm_interconnect_0:mem_master_avalon_master_burstcount
	wire         pcie_ip_bar1_0_waitrequest;                         // mm_interconnect_0:pcie_ip_bar1_0_waitrequest -> pcie_ip:bar1_0_waitrequest
	wire  [63:0] pcie_ip_bar1_0_readdata;                            // mm_interconnect_0:pcie_ip_bar1_0_readdata -> pcie_ip:bar1_0_readdata
	wire  [31:0] pcie_ip_bar1_0_address;                             // pcie_ip:bar1_0_address -> mm_interconnect_0:pcie_ip_bar1_0_address
	wire         pcie_ip_bar1_0_read;                                // pcie_ip:bar1_0_read -> mm_interconnect_0:pcie_ip_bar1_0_read
	wire   [7:0] pcie_ip_bar1_0_byteenable;                          // pcie_ip:bar1_0_byteenable -> mm_interconnect_0:pcie_ip_bar1_0_byteenable
	wire         pcie_ip_bar1_0_readdatavalid;                       // mm_interconnect_0:pcie_ip_bar1_0_readdatavalid -> pcie_ip:bar1_0_readdatavalid
	wire         pcie_ip_bar1_0_write;                               // pcie_ip:bar1_0_write -> mm_interconnect_0:pcie_ip_bar1_0_write
	wire  [63:0] pcie_ip_bar1_0_writedata;                           // pcie_ip:bar1_0_writedata -> mm_interconnect_0:pcie_ip_bar1_0_writedata
	wire   [6:0] pcie_ip_bar1_0_burstcount;                          // pcie_ip:bar1_0_burstcount -> mm_interconnect_0:pcie_ip_bar1_0_burstcount
	wire  [63:0] sgdma_m_read_readdata;                              // mm_interconnect_0:sgdma_m_read_readdata -> sgdma:m_read_readdata
	wire         sgdma_m_read_waitrequest;                           // mm_interconnect_0:sgdma_m_read_waitrequest -> sgdma:m_read_waitrequest
	wire  [31:0] sgdma_m_read_address;                               // sgdma:m_read_address -> mm_interconnect_0:sgdma_m_read_address
	wire         sgdma_m_read_read;                                  // sgdma:m_read_read -> mm_interconnect_0:sgdma_m_read_read
	wire         sgdma_m_read_readdatavalid;                         // mm_interconnect_0:sgdma_m_read_readdatavalid -> sgdma:m_read_readdatavalid
	wire         sgdma_m_write_waitrequest;                          // mm_interconnect_0:sgdma_m_write_waitrequest -> sgdma:m_write_waitrequest
	wire  [31:0] sgdma_m_write_address;                              // sgdma:m_write_address -> mm_interconnect_0:sgdma_m_write_address
	wire   [7:0] sgdma_m_write_byteenable;                           // sgdma:m_write_byteenable -> mm_interconnect_0:sgdma_m_write_byteenable
	wire         sgdma_m_write_write;                                // sgdma:m_write_write -> mm_interconnect_0:sgdma_m_write_write
	wire  [63:0] sgdma_m_write_writedata;                            // sgdma:m_write_writedata -> mm_interconnect_0:sgdma_m_write_writedata
	wire  [31:0] sgdma_descriptor_read_readdata;                     // mm_interconnect_0:sgdma_descriptor_read_readdata -> sgdma:descriptor_read_readdata
	wire         sgdma_descriptor_read_waitrequest;                  // mm_interconnect_0:sgdma_descriptor_read_waitrequest -> sgdma:descriptor_read_waitrequest
	wire  [31:0] sgdma_descriptor_read_address;                      // sgdma:descriptor_read_address -> mm_interconnect_0:sgdma_descriptor_read_address
	wire         sgdma_descriptor_read_read;                         // sgdma:descriptor_read_read -> mm_interconnect_0:sgdma_descriptor_read_read
	wire         sgdma_descriptor_read_readdatavalid;                // mm_interconnect_0:sgdma_descriptor_read_readdatavalid -> sgdma:descriptor_read_readdatavalid
	wire         sgdma_descriptor_write_waitrequest;                 // mm_interconnect_0:sgdma_descriptor_write_waitrequest -> sgdma:descriptor_write_waitrequest
	wire  [31:0] sgdma_descriptor_write_address;                     // sgdma:descriptor_write_address -> mm_interconnect_0:sgdma_descriptor_write_address
	wire         sgdma_descriptor_write_write;                       // sgdma:descriptor_write_write -> mm_interconnect_0:sgdma_descriptor_write_write
	wire  [31:0] sgdma_descriptor_write_writedata;                   // sgdma:descriptor_write_writedata -> mm_interconnect_0:sgdma_descriptor_write_writedata
	wire         mm_interconnect_0_onchip_memory_s1_chipselect;      // mm_interconnect_0:onchip_memory_s1_chipselect -> onchip_memory:chipselect
	wire  [63:0] mm_interconnect_0_onchip_memory_s1_readdata;        // onchip_memory:readdata -> mm_interconnect_0:onchip_memory_s1_readdata
	wire  [13:0] mm_interconnect_0_onchip_memory_s1_address;         // mm_interconnect_0:onchip_memory_s1_address -> onchip_memory:address
	wire   [7:0] mm_interconnect_0_onchip_memory_s1_byteenable;      // mm_interconnect_0:onchip_memory_s1_byteenable -> onchip_memory:byteenable
	wire         mm_interconnect_0_onchip_memory_s1_write;           // mm_interconnect_0:onchip_memory_s1_write -> onchip_memory:write
	wire  [63:0] mm_interconnect_0_onchip_memory_s1_writedata;       // mm_interconnect_0:onchip_memory_s1_writedata -> onchip_memory:writedata
	wire         mm_interconnect_0_onchip_memory_s1_clken;           // mm_interconnect_0:onchip_memory_s1_clken -> onchip_memory:clken
	wire         mm_interconnect_0_sram0_s1_chipselect;              // mm_interconnect_0:sram0_s1_chipselect -> sram0:az_cs
	wire  [31:0] mm_interconnect_0_sram0_s1_readdata;                // sram0:za_data -> mm_interconnect_0:sram0_s1_readdata
	wire         mm_interconnect_0_sram0_s1_waitrequest;             // sram0:za_waitrequest -> mm_interconnect_0:sram0_s1_waitrequest
	wire  [24:0] mm_interconnect_0_sram0_s1_address;                 // mm_interconnect_0:sram0_s1_address -> sram0:az_addr
	wire         mm_interconnect_0_sram0_s1_read;                    // mm_interconnect_0:sram0_s1_read -> sram0:az_rd_n
	wire   [3:0] mm_interconnect_0_sram0_s1_byteenable;              // mm_interconnect_0:sram0_s1_byteenable -> sram0:az_be_n
	wire         mm_interconnect_0_sram0_s1_readdatavalid;           // sram0:za_valid -> mm_interconnect_0:sram0_s1_readdatavalid
	wire         mm_interconnect_0_sram0_s1_write;                   // mm_interconnect_0:sram0_s1_write -> sram0:az_wr_n
	wire  [31:0] mm_interconnect_0_sram0_s1_writedata;               // mm_interconnect_0:sram0_s1_writedata -> sram0:az_data
	wire         mm_interconnect_0_pcie_ip_txs_chipselect;           // mm_interconnect_0:pcie_ip_txs_chipselect -> pcie_ip:txs_chipselect
	wire  [63:0] mm_interconnect_0_pcie_ip_txs_readdata;             // pcie_ip:txs_readdata -> mm_interconnect_0:pcie_ip_txs_readdata
	wire         mm_interconnect_0_pcie_ip_txs_waitrequest;          // pcie_ip:txs_waitrequest -> mm_interconnect_0:pcie_ip_txs_waitrequest
	wire  [30:0] mm_interconnect_0_pcie_ip_txs_address;              // mm_interconnect_0:pcie_ip_txs_address -> pcie_ip:txs_address
	wire         mm_interconnect_0_pcie_ip_txs_read;                 // mm_interconnect_0:pcie_ip_txs_read -> pcie_ip:txs_read
	wire   [7:0] mm_interconnect_0_pcie_ip_txs_byteenable;           // mm_interconnect_0:pcie_ip_txs_byteenable -> pcie_ip:txs_byteenable
	wire         mm_interconnect_0_pcie_ip_txs_readdatavalid;        // pcie_ip:txs_readdatavalid -> mm_interconnect_0:pcie_ip_txs_readdatavalid
	wire         mm_interconnect_0_pcie_ip_txs_write;                // mm_interconnect_0:pcie_ip_txs_write -> pcie_ip:txs_write
	wire  [63:0] mm_interconnect_0_pcie_ip_txs_writedata;            // mm_interconnect_0:pcie_ip_txs_writedata -> pcie_ip:txs_writedata
	wire   [6:0] mm_interconnect_0_pcie_ip_txs_burstcount;           // mm_interconnect_0:pcie_ip_txs_burstcount -> pcie_ip:txs_burstcount
	wire  [31:0] mm_interconnect_0_ssram0_uas_readdata;              // ssram0:uas_readdata -> mm_interconnect_0:ssram0_uas_readdata
	wire         mm_interconnect_0_ssram0_uas_waitrequest;           // ssram0:uas_waitrequest -> mm_interconnect_0:ssram0_uas_waitrequest
	wire         mm_interconnect_0_ssram0_uas_debugaccess;           // mm_interconnect_0:ssram0_uas_debugaccess -> ssram0:uas_debugaccess
	wire  [21:0] mm_interconnect_0_ssram0_uas_address;               // mm_interconnect_0:ssram0_uas_address -> ssram0:uas_address
	wire         mm_interconnect_0_ssram0_uas_read;                  // mm_interconnect_0:ssram0_uas_read -> ssram0:uas_read
	wire   [3:0] mm_interconnect_0_ssram0_uas_byteenable;            // mm_interconnect_0:ssram0_uas_byteenable -> ssram0:uas_byteenable
	wire         mm_interconnect_0_ssram0_uas_readdatavalid;         // ssram0:uas_readdatavalid -> mm_interconnect_0:ssram0_uas_readdatavalid
	wire         mm_interconnect_0_ssram0_uas_lock;                  // mm_interconnect_0:ssram0_uas_lock -> ssram0:uas_lock
	wire         mm_interconnect_0_ssram0_uas_write;                 // mm_interconnect_0:ssram0_uas_write -> ssram0:uas_write
	wire  [31:0] mm_interconnect_0_ssram0_uas_writedata;             // mm_interconnect_0:ssram0_uas_writedata -> ssram0:uas_writedata
	wire   [2:0] mm_interconnect_0_ssram0_uas_burstcount;            // mm_interconnect_0:ssram0_uas_burstcount -> ssram0:uas_burstcount
	wire  [31:0] mm_interconnect_0_ssram1_uas_readdata;              // ssram1:uas_readdata -> mm_interconnect_0:ssram1_uas_readdata
	wire         mm_interconnect_0_ssram1_uas_waitrequest;           // ssram1:uas_waitrequest -> mm_interconnect_0:ssram1_uas_waitrequest
	wire         mm_interconnect_0_ssram1_uas_debugaccess;           // mm_interconnect_0:ssram1_uas_debugaccess -> ssram1:uas_debugaccess
	wire  [21:0] mm_interconnect_0_ssram1_uas_address;               // mm_interconnect_0:ssram1_uas_address -> ssram1:uas_address
	wire         mm_interconnect_0_ssram1_uas_read;                  // mm_interconnect_0:ssram1_uas_read -> ssram1:uas_read
	wire   [3:0] mm_interconnect_0_ssram1_uas_byteenable;            // mm_interconnect_0:ssram1_uas_byteenable -> ssram1:uas_byteenable
	wire         mm_interconnect_0_ssram1_uas_readdatavalid;         // ssram1:uas_readdatavalid -> mm_interconnect_0:ssram1_uas_readdatavalid
	wire         mm_interconnect_0_ssram1_uas_lock;                  // mm_interconnect_0:ssram1_uas_lock -> ssram1:uas_lock
	wire         mm_interconnect_0_ssram1_uas_write;                 // mm_interconnect_0:ssram1_uas_write -> ssram1:uas_write
	wire  [31:0] mm_interconnect_0_ssram1_uas_writedata;             // mm_interconnect_0:ssram1_uas_writedata -> ssram1:uas_writedata
	wire   [2:0] mm_interconnect_0_ssram1_uas_burstcount;            // mm_interconnect_0:ssram1_uas_burstcount -> ssram1:uas_burstcount
	wire         mm_interconnect_0_led_s1_chipselect;                // mm_interconnect_0:led_s1_chipselect -> led:chipselect
	wire  [31:0] mm_interconnect_0_led_s1_readdata;                  // led:readdata -> mm_interconnect_0:led_s1_readdata
	wire   [1:0] mm_interconnect_0_led_s1_address;                   // mm_interconnect_0:led_s1_address -> led:address
	wire         mm_interconnect_0_led_s1_write;                     // mm_interconnect_0:led_s1_write -> led:write_n
	wire  [31:0] mm_interconnect_0_led_s1_writedata;                 // mm_interconnect_0:led_s1_writedata -> led:writedata
	wire         mm_interconnect_0_button_s1_chipselect;             // mm_interconnect_0:button_s1_chipselect -> button:chipselect
	wire  [31:0] mm_interconnect_0_button_s1_readdata;               // button:readdata -> mm_interconnect_0:button_s1_readdata
	wire   [1:0] mm_interconnect_0_button_s1_address;                // mm_interconnect_0:button_s1_address -> button:address
	wire         mm_interconnect_0_button_s1_write;                  // mm_interconnect_0:button_s1_write -> button:write_n
	wire  [31:0] mm_interconnect_0_button_s1_writedata;              // mm_interconnect_0:button_s1_writedata -> button:writedata
	wire         mm_interconnect_0_pio_size_s1_chipselect;           // mm_interconnect_0:pio_size_s1_chipselect -> pio_size:chipselect
	wire  [31:0] mm_interconnect_0_pio_size_s1_readdata;             // pio_size:readdata -> mm_interconnect_0:pio_size_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_size_s1_address;              // mm_interconnect_0:pio_size_s1_address -> pio_size:address
	wire         mm_interconnect_0_pio_size_s1_write;                // mm_interconnect_0:pio_size_s1_write -> pio_size:write_n
	wire  [31:0] mm_interconnect_0_pio_size_s1_writedata;            // mm_interconnect_0:pio_size_s1_writedata -> pio_size:writedata
	wire         mm_interconnect_0_chip_sel_s1_chipselect;           // mm_interconnect_0:chip_sel_s1_chipselect -> chip_sel:chipselect
	wire  [31:0] mm_interconnect_0_chip_sel_s1_readdata;             // chip_sel:readdata -> mm_interconnect_0:chip_sel_s1_readdata
	wire   [1:0] mm_interconnect_0_chip_sel_s1_address;              // mm_interconnect_0:chip_sel_s1_address -> chip_sel:address
	wire         mm_interconnect_0_chip_sel_s1_write;                // mm_interconnect_0:chip_sel_s1_write -> chip_sel:write_n
	wire  [31:0] mm_interconnect_0_chip_sel_s1_writedata;            // mm_interconnect_0:chip_sel_s1_writedata -> chip_sel:writedata
	wire  [31:0] mm_interconnect_0_width_s1_readdata;                // width:readdata -> mm_interconnect_0:width_s1_readdata
	wire   [1:0] mm_interconnect_0_width_s1_address;                 // mm_interconnect_0:width_s1_address -> width:address
	wire  [31:0] mm_interconnect_0_height_s1_readdata;               // height:readdata -> mm_interconnect_0:height_s1_readdata
	wire   [1:0] mm_interconnect_0_height_s1_address;                // mm_interconnect_0:height_s1_address -> height:address
	wire         pcie_ip_bar2_waitrequest;                           // mm_interconnect_1:pcie_ip_bar2_waitrequest -> pcie_ip:bar2_waitrequest
	wire  [63:0] pcie_ip_bar2_readdata;                              // mm_interconnect_1:pcie_ip_bar2_readdata -> pcie_ip:bar2_readdata
	wire  [31:0] pcie_ip_bar2_address;                               // pcie_ip:bar2_address -> mm_interconnect_1:pcie_ip_bar2_address
	wire         pcie_ip_bar2_read;                                  // pcie_ip:bar2_read -> mm_interconnect_1:pcie_ip_bar2_read
	wire   [7:0] pcie_ip_bar2_byteenable;                            // pcie_ip:bar2_byteenable -> mm_interconnect_1:pcie_ip_bar2_byteenable
	wire         pcie_ip_bar2_readdatavalid;                         // mm_interconnect_1:pcie_ip_bar2_readdatavalid -> pcie_ip:bar2_readdatavalid
	wire         pcie_ip_bar2_write;                                 // pcie_ip:bar2_write -> mm_interconnect_1:pcie_ip_bar2_write
	wire  [63:0] pcie_ip_bar2_writedata;                             // pcie_ip:bar2_writedata -> mm_interconnect_1:pcie_ip_bar2_writedata
	wire   [6:0] pcie_ip_bar2_burstcount;                            // pcie_ip:bar2_burstcount -> mm_interconnect_1:pcie_ip_bar2_burstcount
	wire         mm_interconnect_1_pcie_ip_cra_chipselect;           // mm_interconnect_1:pcie_ip_cra_chipselect -> pcie_ip:cra_chipselect
	wire  [31:0] mm_interconnect_1_pcie_ip_cra_readdata;             // pcie_ip:cra_readdata -> mm_interconnect_1:pcie_ip_cra_readdata
	wire         mm_interconnect_1_pcie_ip_cra_waitrequest;          // pcie_ip:cra_waitrequest -> mm_interconnect_1:pcie_ip_cra_waitrequest
	wire  [11:0] mm_interconnect_1_pcie_ip_cra_address;              // mm_interconnect_1:pcie_ip_cra_address -> pcie_ip:cra_address
	wire         mm_interconnect_1_pcie_ip_cra_read;                 // mm_interconnect_1:pcie_ip_cra_read -> pcie_ip:cra_read
	wire   [3:0] mm_interconnect_1_pcie_ip_cra_byteenable;           // mm_interconnect_1:pcie_ip_cra_byteenable -> pcie_ip:cra_byteenable
	wire         mm_interconnect_1_pcie_ip_cra_write;                // mm_interconnect_1:pcie_ip_cra_write -> pcie_ip:cra_write
	wire  [31:0] mm_interconnect_1_pcie_ip_cra_writedata;            // mm_interconnect_1:pcie_ip_cra_writedata -> pcie_ip:cra_writedata
	wire         mm_interconnect_1_sgdma_csr_chipselect;             // mm_interconnect_1:sgdma_csr_chipselect -> sgdma:csr_chipselect
	wire  [31:0] mm_interconnect_1_sgdma_csr_readdata;               // sgdma:csr_readdata -> mm_interconnect_1:sgdma_csr_readdata
	wire   [3:0] mm_interconnect_1_sgdma_csr_address;                // mm_interconnect_1:sgdma_csr_address -> sgdma:csr_address
	wire         mm_interconnect_1_sgdma_csr_read;                   // mm_interconnect_1:sgdma_csr_read -> sgdma:csr_read
	wire         mm_interconnect_1_sgdma_csr_write;                  // mm_interconnect_1:sgdma_csr_write -> sgdma:csr_write
	wire  [31:0] mm_interconnect_1_sgdma_csr_writedata;              // mm_interconnect_1:sgdma_csr_writedata -> sgdma:csr_writedata
	wire         irq_mapper_receiver0_irq;                           // sgdma:csr_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                           // button:irq -> irq_mapper:receiver1_irq
	wire  [15:0] pcie_ip_rxm_irq_irq;                                // irq_mapper:sender_irq -> pcie_ip:rxm_irq_irq
	wire         rst_controller_reset_out_reset;                     // rst_controller:reset_out -> altpll_0:reset
	wire         pcie_ip_pcie_core_reset_reset;                      // pcie_ip:pcie_core_reset_reset_n -> [rst_controller:reset_in1, rst_controller_001:reset_in1, rst_controller_002:reset_in1, rst_controller_003:reset_in0]
	wire         rst_controller_001_reset_out_reset;                 // rst_controller_001:reset_out -> [button:reset_n, chip_sel:reset_n, height:reset_n, led:reset_n, mem_master:reset, mm_interconnect_0:mem_master_clock_reset_reset_reset_bridge_in_reset_reset, mm_interconnect_1:sgdma_reset_reset_bridge_in_reset_reset, onchip_memory:reset, onchip_memory:reset2, pio_size:reset_n, rst_controller_001_reset_out_reset:in, rst_translator:in_reset, sgdma:system_reset_n, ssram0:reset_reset, ssram1:reset_reset, tristate_conduit_bridge_0:reset, tristate_conduit_pin_sharer_0:reset_reset, width:reset_n]
	wire         rst_controller_001_reset_out_reset_req;             // rst_controller_001:reset_req -> [onchip_memory:reset_req, onchip_memory:reset_req2, rst_translator:reset_req_in]
	wire         rst_controller_002_reset_out_reset;                 // rst_controller_002:reset_out -> [mm_interconnect_0:sram0_reset_reset_bridge_in_reset_reset, sram0:reset_n]
	wire         rst_controller_003_reset_out_reset;                 // rst_controller_003:reset_out -> [irq_mapper:reset, mm_interconnect_0:pcie_ip_bar1_0_translator_reset_reset_bridge_in_reset_reset, mm_interconnect_1:pcie_ip_bar2_translator_reset_reset_bridge_in_reset_reset]

	de2i_150_qsys_altpll_0 altpll_0 (
		.clk       (clk_clk),                        //       inclk_interface.clk
		.reset     (rst_controller_reset_out_reset), // inclk_interface_reset.reset
		.read      (),                               //             pll_slave.read
		.write     (),                               //                      .write
		.address   (),                               //                      .address
		.readdata  (),                               //                      .readdata
		.writedata (),                               //                      .writedata
		.c0        (altpll_sdram_clk),               //                    c0.clk
		.c1        (altpll_0_c1_clk),                //                    c1.clk
		.areset    (),                               //        areset_conduit.export
		.locked    (),                               //        locked_conduit.export
		.phasedone ()                                //     phasedone_conduit.export
	);

	de2i_150_qsys_button button (
		.clk        (pcie_clk_clk),                           //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),    //               reset.reset_n
		.address    (mm_interconnect_0_button_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_button_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_button_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_button_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_button_s1_readdata),   //                    .readdata
		.in_port    (button_external_connection_export),      // external_connection.export
		.irq        (irq_mapper_receiver1_irq)                //                 irq.irq
	);

	de2i_150_qsys_chip_sel chip_sel (
		.clk        (pcie_clk_clk),                             //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_chip_sel_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_chip_sel_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_chip_sel_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_chip_sel_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_chip_sel_s1_readdata),   //                    .readdata
		.out_port   (chip_sel_export)                           // external_connection.export
	);

	de2i_150_qsys_height height (
		.clk      (pcie_clk_clk),                         //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),  //               reset.reset_n
		.address  (mm_interconnect_0_height_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_height_s1_readdata), //                    .readdata
		.in_port  (height_external_connection_export)     // external_connection.export
	);

	de2i_150_qsys_led led (
		.clk        (pcie_clk_clk),                        //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset), //               reset.reset_n
		.address    (mm_interconnect_0_led_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_led_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_led_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_led_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_led_s1_readdata),   //                    .readdata
		.out_port   (led_external_connection_export)       // external_connection.export
	);

	custom_master #(
		.MASTER_DIRECTION    (0),
		.DATA_WIDTH          (32),
		.ADDRESS_WIDTH       (32),
		.BURST_CAPABLE       (1),
		.MAXIMUM_BURST_COUNT (128),
		.BURST_COUNT_WIDTH   (8),
		.FIFO_DEPTH          (256),
		.FIFO_DEPTH_LOG2     (8),
		.MEMORY_BASED_FIFO   (1)
	) mem_master (
		.clk                     (pcie_clk_clk),                           //       clock_reset.clk
		.reset                   (rst_controller_001_reset_out_reset),     // clock_reset_reset.reset
		.master_address          (mem_master_avalon_master_address),       //     avalon_master.address
		.master_read             (mem_master_avalon_master_read),          //                  .read
		.master_byteenable       (mem_master_avalon_master_byteenable),    //                  .byteenable
		.master_readdata         (mem_master_avalon_master_readdata),      //                  .readdata
		.master_readdatavalid    (mem_master_avalon_master_readdatavalid), //                  .readdatavalid
		.master_burstcount       (mem_master_avalon_master_burstcount),    //                  .burstcount
		.master_waitrequest      (mem_master_avalon_master_waitrequest),   //                  .waitrequest
		.control_fixed_location  (mem_master_control_fixed_location),      //           control.export
		.control_read_base       (mem_master_control_read_base),           //                  .export
		.control_read_length     (mem_master_control_read_length),         //                  .export
		.control_go              (mem_master_control_go),                  //                  .export
		.control_done            (mem_master_control_done),                //                  .export
		.control_early_done      (mem_master_control_early_done),          //                  .export
		.user_read_buffer        (mem_master_user_read_buffer),            //              user.export
		.user_buffer_output_data (mem_master_user_buffer_output_data),     //                  .export
		.user_data_available     (mem_master_user_data_available),         //                  .export
		.master_write            (),                                       //       (terminated)
		.master_writedata        (),                                       //       (terminated)
		.control_write_base      (32'b00000000000000000000000000000000),   //       (terminated)
		.control_write_length    (32'b00000000000000000000000000000000),   //       (terminated)
		.user_write_buffer       (1'b0),                                   //       (terminated)
		.user_buffer_input_data  (32'b00000000000000000000000000000000),   //       (terminated)
		.user_buffer_full        ()                                        //       (terminated)
	);

	de2i_150_qsys_onchip_memory onchip_memory (
		.clk         (pcie_clk_clk),                                  //   clk1.clk
		.address     (mm_interconnect_0_onchip_memory_s1_address),    //     s1.address
		.clken       (mm_interconnect_0_onchip_memory_s1_clken),      //       .clken
		.chipselect  (mm_interconnect_0_onchip_memory_s1_chipselect), //       .chipselect
		.write       (mm_interconnect_0_onchip_memory_s1_write),      //       .write
		.readdata    (mm_interconnect_0_onchip_memory_s1_readdata),   //       .readdata
		.writedata   (mm_interconnect_0_onchip_memory_s1_writedata),  //       .writedata
		.byteenable  (mm_interconnect_0_onchip_memory_s1_byteenable), //       .byteenable
		.reset       (rst_controller_001_reset_out_reset),            // reset1.reset
		.reset_req   (rst_controller_001_reset_out_reset_req),        //       .reset_req
		.address2    (),                                              //     s2.address
		.chipselect2 (),                                              //       .chipselect
		.clken2      (),                                              //       .clken
		.write2      (),                                              //       .write
		.readdata2   (),                                              //       .readdata
		.writedata2  (),                                              //       .writedata
		.byteenable2 (),                                              //       .byteenable
		.clk2        (pcie_clk_clk),                                  //   clk2.clk
		.reset2      (rst_controller_001_reset_out_reset),            // reset2.reset
		.reset_req2  (rst_controller_001_reset_out_reset_req)         //       .reset_req
	);

	de2i_150_qsys_pcie_ip #(
		.p_pcie_hip_type                     ("2"),
		.lane_mask                           (8'b11111110),
		.max_link_width                      (1),
		.millisecond_cycle_count             ("125000"),
		.enable_gen2_core                    ("false"),
		.gen2_lane_rate_mode                 ("false"),
		.no_soft_reset                       ("false"),
		.core_clk_divider                    (2),
		.enable_ch0_pclk_out                 ("true"),
		.core_clk_source                     ("pclk"),
		.CB_P2A_AVALON_ADDR_B0               (0),
		.bar0_size_mask                      (28),
		.bar0_io_space                       ("false"),
		.bar0_64bit_mem_space                ("true"),
		.bar0_prefetchable                   ("true"),
		.CB_P2A_AVALON_ADDR_B1               (0),
		.bar1_size_mask                      (0),
		.bar1_io_space                       ("false"),
		.bar1_64bit_mem_space                ("true"),
		.bar1_prefetchable                   ("false"),
		.CB_P2A_AVALON_ADDR_B2               (0),
		.bar2_size_mask                      (15),
		.bar2_io_space                       ("false"),
		.bar2_64bit_mem_space                ("false"),
		.bar2_prefetchable                   ("false"),
		.CB_P2A_AVALON_ADDR_B3               (0),
		.bar3_size_mask                      (0),
		.bar3_io_space                       ("false"),
		.bar3_64bit_mem_space                ("false"),
		.bar3_prefetchable                   ("false"),
		.CB_P2A_AVALON_ADDR_B4               (0),
		.bar4_size_mask                      (0),
		.bar4_io_space                       ("false"),
		.bar4_64bit_mem_space                ("false"),
		.bar4_prefetchable                   ("false"),
		.CB_P2A_AVALON_ADDR_B5               (0),
		.bar5_size_mask                      (0),
		.bar5_io_space                       ("false"),
		.bar5_64bit_mem_space                ("false"),
		.bar5_prefetchable                   ("false"),
		.vendor_id                           (4466),
		.device_id                           (57345),
		.revision_id                         (1),
		.class_code                          (0),
		.subsystem_vendor_id                 (4466),
		.subsystem_device_id                 (4),
		.port_link_number                    (1),
		.msi_function_count                  (0),
		.enable_msi_64bit_addressing         ("true"),
		.enable_function_msix_support        ("false"),
		.eie_before_nfts_count               (4),
		.enable_completion_timeout_disable   ("false"),
		.completion_timeout                  ("NONE"),
		.enable_adapter_half_rate_mode       ("false"),
		.msix_pba_bir                        (0),
		.msix_pba_offset                     (0),
		.msix_table_bir                      (0),
		.msix_table_offset                   (0),
		.msix_table_size                     (0),
		.use_crc_forwarding                  ("false"),
		.surprise_down_error_support         ("false"),
		.dll_active_report_support           ("false"),
		.bar_io_window_size                  ("32BIT"),
		.bar_prefetchable                    (32),
		.hot_plug_support                    (7'b0000000),
		.no_command_completed                ("true"),
		.slot_power_limit                    (0),
		.slot_power_scale                    (0),
		.slot_number                         (0),
		.enable_slot_register                ("false"),
		.advanced_errors                     ("false"),
		.enable_ecrc_check                   ("false"),
		.enable_ecrc_gen                     ("false"),
		.max_payload_size                    (0),
		.retry_buffer_last_active_address    (255),
		.credit_buffer_allocation_aux        ("ABSOLUTE"),
		.vc0_rx_flow_ctrl_posted_header      (28),
		.vc0_rx_flow_ctrl_posted_data        (198),
		.vc0_rx_flow_ctrl_nonposted_header   (30),
		.vc0_rx_flow_ctrl_nonposted_data     (0),
		.vc0_rx_flow_ctrl_compl_header       (48),
		.vc0_rx_flow_ctrl_compl_data         (256),
		.RX_BUF                              (9),
		.RH_NUM                              (7),
		.G_TAG_NUM0                          (32),
		.endpoint_l0_latency                 (0),
		.endpoint_l1_latency                 (0),
		.enable_l1_aspm                      ("false"),
		.l01_entry_latency                   (31),
		.diffclock_nfts_count                (255),
		.sameclock_nfts_count                (255),
		.l1_exit_latency_sameclock           (7),
		.l1_exit_latency_diffclock           (7),
		.l0_exit_latency_sameclock           (7),
		.l0_exit_latency_diffclock           (7),
		.gen2_diffclock_nfts_count           (255),
		.gen2_sameclock_nfts_count           (255),
		.CG_COMMON_CLOCK_MODE                (1),
		.CB_PCIE_MODE                        (0),
		.AST_LITE                            (0),
		.CB_PCIE_RX_LITE                     (0),
		.CG_RXM_IRQ_NUM                      (16),
		.CG_AVALON_S_ADDR_WIDTH              (20),
		.bypass_tl                           ("false"),
		.CG_IMPL_CRA_AV_SLAVE_PORT           (1),
		.CG_NO_CPL_REORDERING                (0),
		.CG_ENABLE_A2P_INTERRUPT             (0),
		.p_user_msi_enable                   (0),
		.CG_IRQ_BIT_ENA                      (65535),
		.CB_A2P_ADDR_MAP_IS_FIXED            (1),
		.CB_A2P_ADDR_MAP_NUM_ENTRIES         (1),
		.CB_A2P_ADDR_MAP_PASS_THRU_BITS      (31),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_0_HIGH  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_0_LOW   (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_1_HIGH  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_1_LOW   (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_2_HIGH  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_2_LOW   (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_3_HIGH  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_3_LOW   (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_4_HIGH  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_4_LOW   (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_5_HIGH  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_5_LOW   (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_6_HIGH  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_6_LOW   (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_7_HIGH  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_7_LOW   (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_8_HIGH  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_8_LOW   (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_9_HIGH  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_9_LOW   (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_10_HIGH (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_10_LOW  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_11_HIGH (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_11_LOW  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_12_HIGH (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_12_LOW  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_13_HIGH (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_13_LOW  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_14_HIGH (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_14_LOW  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_15_HIGH (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_15_LOW  (32'b00000000000000000000000000000000),
		.RXM_DATA_WIDTH                      (64),
		.RXM_BEN_WIDTH                       (8),
		.TL_SELECTION                        (1),
		.pcie_mode                           ("SHARED_MODE"),
		.single_rx_detect                    (1),
		.enable_coreclk_out_half_rate        ("false"),
		.low_priority_vc                     (0),
		.link_width                          (1),
		.cyclone4                            (1)
	) pcie_ip (
		.pcie_core_clk_clk                  (pcie_clk_clk),                                //      pcie_core_clk.clk
		.pcie_core_reset_reset_n            (pcie_ip_pcie_core_reset_reset),               //    pcie_core_reset.reset_n
		.cal_blk_clk_clk                    (clk_clk),                                     //        cal_blk_clk.clk
		.txs_address                        (mm_interconnect_0_pcie_ip_txs_address),       //                txs.address
		.txs_chipselect                     (mm_interconnect_0_pcie_ip_txs_chipselect),    //                   .chipselect
		.txs_byteenable                     (mm_interconnect_0_pcie_ip_txs_byteenable),    //                   .byteenable
		.txs_readdata                       (mm_interconnect_0_pcie_ip_txs_readdata),      //                   .readdata
		.txs_writedata                      (mm_interconnect_0_pcie_ip_txs_writedata),     //                   .writedata
		.txs_read                           (mm_interconnect_0_pcie_ip_txs_read),          //                   .read
		.txs_write                          (mm_interconnect_0_pcie_ip_txs_write),         //                   .write
		.txs_burstcount                     (mm_interconnect_0_pcie_ip_txs_burstcount),    //                   .burstcount
		.txs_readdatavalid                  (mm_interconnect_0_pcie_ip_txs_readdatavalid), //                   .readdatavalid
		.txs_waitrequest                    (mm_interconnect_0_pcie_ip_txs_waitrequest),   //                   .waitrequest
		.refclk_export                      (pcie_ip_refclk_export),                       //             refclk.export
		.test_in_test_in                    (pcie_ip_test_in_test_in),                     //            test_in.test_in
		.pcie_rstn_export                   (pcie_ip_pcie_rstn_export),                    //          pcie_rstn.export
		.clocks_sim_clk250_export           (pcie_ip_clocks_sim_clk250_export),            //         clocks_sim.clk250_export
		.clocks_sim_clk500_export           (pcie_ip_clocks_sim_clk500_export),            //                   .clk500_export
		.clocks_sim_clk125_export           (pcie_ip_clocks_sim_clk125_export),            //                   .clk125_export
		.reconfig_busy_busy_altgxb_reconfig (pcie_ip_reconfig_busy_busy_altgxb_reconfig),  //      reconfig_busy.busy_altgxb_reconfig
		.pipe_ext_pipe_mode                 (pcie_ip_pipe_ext_pipe_mode),                  //           pipe_ext.pipe_mode
		.pipe_ext_phystatus_ext             (pcie_ip_pipe_ext_phystatus_ext),              //                   .phystatus_ext
		.pipe_ext_rate_ext                  (pcie_ip_pipe_ext_rate_ext),                   //                   .rate_ext
		.pipe_ext_powerdown_ext             (pcie_ip_pipe_ext_powerdown_ext),              //                   .powerdown_ext
		.pipe_ext_txdetectrx_ext            (pcie_ip_pipe_ext_txdetectrx_ext),             //                   .txdetectrx_ext
		.pipe_ext_rxelecidle0_ext           (pcie_ip_pipe_ext_rxelecidle0_ext),            //                   .rxelecidle0_ext
		.pipe_ext_rxdata0_ext               (pcie_ip_pipe_ext_rxdata0_ext),                //                   .rxdata0_ext
		.pipe_ext_rxstatus0_ext             (pcie_ip_pipe_ext_rxstatus0_ext),              //                   .rxstatus0_ext
		.pipe_ext_rxvalid0_ext              (pcie_ip_pipe_ext_rxvalid0_ext),               //                   .rxvalid0_ext
		.pipe_ext_rxdatak0_ext              (pcie_ip_pipe_ext_rxdatak0_ext),               //                   .rxdatak0_ext
		.pipe_ext_txdata0_ext               (pcie_ip_pipe_ext_txdata0_ext),                //                   .txdata0_ext
		.pipe_ext_txdatak0_ext              (pcie_ip_pipe_ext_txdatak0_ext),               //                   .txdatak0_ext
		.pipe_ext_rxpolarity0_ext           (pcie_ip_pipe_ext_rxpolarity0_ext),            //                   .rxpolarity0_ext
		.pipe_ext_txcompl0_ext              (pcie_ip_pipe_ext_txcompl0_ext),               //                   .txcompl0_ext
		.pipe_ext_txelecidle0_ext           (pcie_ip_pipe_ext_txelecidle0_ext),            //                   .txelecidle0_ext
		.powerdown_pll_powerdown            (),                                            //          powerdown.pll_powerdown
		.powerdown_gxb_powerdown            (),                                            //                   .gxb_powerdown
		.bar1_0_address                     (pcie_ip_bar1_0_address),                      //             bar1_0.address
		.bar1_0_read                        (pcie_ip_bar1_0_read),                         //                   .read
		.bar1_0_waitrequest                 (pcie_ip_bar1_0_waitrequest),                  //                   .waitrequest
		.bar1_0_write                       (pcie_ip_bar1_0_write),                        //                   .write
		.bar1_0_readdatavalid               (pcie_ip_bar1_0_readdatavalid),                //                   .readdatavalid
		.bar1_0_readdata                    (pcie_ip_bar1_0_readdata),                     //                   .readdata
		.bar1_0_writedata                   (pcie_ip_bar1_0_writedata),                    //                   .writedata
		.bar1_0_burstcount                  (pcie_ip_bar1_0_burstcount),                   //                   .burstcount
		.bar1_0_byteenable                  (pcie_ip_bar1_0_byteenable),                   //                   .byteenable
		.bar2_address                       (pcie_ip_bar2_address),                        //               bar2.address
		.bar2_read                          (pcie_ip_bar2_read),                           //                   .read
		.bar2_waitrequest                   (pcie_ip_bar2_waitrequest),                    //                   .waitrequest
		.bar2_write                         (pcie_ip_bar2_write),                          //                   .write
		.bar2_readdatavalid                 (pcie_ip_bar2_readdatavalid),                  //                   .readdatavalid
		.bar2_readdata                      (pcie_ip_bar2_readdata),                       //                   .readdata
		.bar2_writedata                     (pcie_ip_bar2_writedata),                      //                   .writedata
		.bar2_burstcount                    (pcie_ip_bar2_burstcount),                     //                   .burstcount
		.bar2_byteenable                    (pcie_ip_bar2_byteenable),                     //                   .byteenable
		.cra_chipselect                     (mm_interconnect_1_pcie_ip_cra_chipselect),    //                cra.chipselect
		.cra_address                        (mm_interconnect_1_pcie_ip_cra_address),       //                   .address
		.cra_byteenable                     (mm_interconnect_1_pcie_ip_cra_byteenable),    //                   .byteenable
		.cra_read                           (mm_interconnect_1_pcie_ip_cra_read),          //                   .read
		.cra_readdata                       (mm_interconnect_1_pcie_ip_cra_readdata),      //                   .readdata
		.cra_write                          (mm_interconnect_1_pcie_ip_cra_write),         //                   .write
		.cra_writedata                      (mm_interconnect_1_pcie_ip_cra_writedata),     //                   .writedata
		.cra_waitrequest                    (mm_interconnect_1_pcie_ip_cra_waitrequest),   //                   .waitrequest
		.cra_irq_irq                        (),                                            //            cra_irq.irq
		.rxm_irq_irq                        (pcie_ip_rxm_irq_irq),                         //            rxm_irq.irq
		.rx_in_rx_datain_0                  (pcie_ip_rx_in_rx_datain_0),                   //              rx_in.rx_datain_0
		.tx_out_tx_dataout_0                (pcie_ip_tx_out_tx_dataout_0),                 //             tx_out.tx_dataout_0
		.reconfig_togxb_data                (pcie_ip_reconfig_togxb_data),                 //     reconfig_togxb.data
		.reconfig_gxbclk_clk                (clk_clk),                                     //    reconfig_gxbclk.clk
		.reconfig_fromgxb_0_data            (pcie_ip_reconfig_fromgxb_0_data),             // reconfig_fromgxb_0.data
		.fixedclk_clk                       (pcie_clk_clk)                                 //           fixedclk.clk
	);

	de2i_150_qsys_pio_size pio_size (
		.clk        (pcie_clk_clk),                             //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_pio_size_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_size_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_size_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_size_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_size_s1_readdata),   //                    .readdata
		.out_port   (pio_size_external_connection_export)       // external_connection.export
	);

	de2i_150_qsys_sgdma sgdma (
		.clk                           (pcie_clk_clk),                           //              clk.clk
		.system_reset_n                (~rst_controller_001_reset_out_reset),    //            reset.reset_n
		.csr_chipselect                (mm_interconnect_1_sgdma_csr_chipselect), //              csr.chipselect
		.csr_address                   (mm_interconnect_1_sgdma_csr_address),    //                 .address
		.csr_read                      (mm_interconnect_1_sgdma_csr_read),       //                 .read
		.csr_write                     (mm_interconnect_1_sgdma_csr_write),      //                 .write
		.csr_writedata                 (mm_interconnect_1_sgdma_csr_writedata),  //                 .writedata
		.csr_readdata                  (mm_interconnect_1_sgdma_csr_readdata),   //                 .readdata
		.descriptor_read_readdata      (sgdma_descriptor_read_readdata),         //  descriptor_read.readdata
		.descriptor_read_readdatavalid (sgdma_descriptor_read_readdatavalid),    //                 .readdatavalid
		.descriptor_read_waitrequest   (sgdma_descriptor_read_waitrequest),      //                 .waitrequest
		.descriptor_read_address       (sgdma_descriptor_read_address),          //                 .address
		.descriptor_read_read          (sgdma_descriptor_read_read),             //                 .read
		.descriptor_write_waitrequest  (sgdma_descriptor_write_waitrequest),     // descriptor_write.waitrequest
		.descriptor_write_address      (sgdma_descriptor_write_address),         //                 .address
		.descriptor_write_write        (sgdma_descriptor_write_write),           //                 .write
		.descriptor_write_writedata    (sgdma_descriptor_write_writedata),       //                 .writedata
		.csr_irq                       (irq_mapper_receiver0_irq),               //          csr_irq.irq
		.m_read_readdata               (sgdma_m_read_readdata),                  //           m_read.readdata
		.m_read_readdatavalid          (sgdma_m_read_readdatavalid),             //                 .readdatavalid
		.m_read_waitrequest            (sgdma_m_read_waitrequest),               //                 .waitrequest
		.m_read_address                (sgdma_m_read_address),                   //                 .address
		.m_read_read                   (sgdma_m_read_read),                      //                 .read
		.m_write_waitrequest           (sgdma_m_write_waitrequest),              //          m_write.waitrequest
		.m_write_address               (sgdma_m_write_address),                  //                 .address
		.m_write_write                 (sgdma_m_write_write),                    //                 .write
		.m_write_writedata             (sgdma_m_write_writedata),                //                 .writedata
		.m_write_byteenable            (sgdma_m_write_byteenable)                //                 .byteenable
	);

	de2i_150_qsys_sram0 sram0 (
		.clk            (altpll_0_c1_clk),                          //   clk.clk
		.reset_n        (~rst_controller_002_reset_out_reset),      // reset.reset_n
		.az_addr        (mm_interconnect_0_sram0_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sram0_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sram0_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sram0_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sram0_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sram0_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sram0_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sram0_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sram0_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_addr),                               //  wire.export
		.zs_ba          (sdram_ba),                                 //      .export
		.zs_cas_n       (sdram_cas_n),                              //      .export
		.zs_cke         (sdram_cke),                                //      .export
		.zs_cs_n        (sdram_cs_n),                               //      .export
		.zs_dq          (sdram_dq),                                 //      .export
		.zs_dqm         (sdram_dqm),                                //      .export
		.zs_ras_n       (sdram_ras_n),                              //      .export
		.zs_we_n        (sdram_we_n)                                //      .export
	);

	de2i_150_qsys_ssram0 #(
		.TCM_ADDRESS_W                  (22),
		.TCM_DATA_W                     (32),
		.TCM_BYTEENABLE_W               (4),
		.TCM_READ_WAIT                  (0),
		.TCM_WRITE_WAIT                 (0),
		.TCM_SETUP_WAIT                 (0),
		.TCM_DATA_HOLD                  (0),
		.TCM_TURNAROUND_TIME            (2),
		.TCM_TIMING_UNITS               (1),
		.TCM_READLATENCY                (4),
		.TCM_SYMBOLS_PER_WORD           (4),
		.USE_READDATA                   (1),
		.USE_WRITEDATA                  (1),
		.USE_READ                       (0),
		.USE_WRITE                      (1),
		.USE_BYTEENABLE                 (1),
		.USE_CHIPSELECT                 (1),
		.USE_LOCK                       (0),
		.USE_ADDRESS                    (1),
		.USE_WAITREQUEST                (0),
		.USE_WRITEBYTEENABLE            (0),
		.USE_OUTPUTENABLE               (1),
		.USE_RESETREQUEST               (0),
		.USE_IRQ                        (0),
		.USE_RESET_OUTPUT               (0),
		.ACTIVE_LOW_READ                (0),
		.ACTIVE_LOW_LOCK                (0),
		.ACTIVE_LOW_WRITE               (1),
		.ACTIVE_LOW_CHIPSELECT          (1),
		.ACTIVE_LOW_BYTEENABLE          (1),
		.ACTIVE_LOW_OUTPUTENABLE        (1),
		.ACTIVE_LOW_WRITEBYTEENABLE     (0),
		.ACTIVE_LOW_WAITREQUEST         (0),
		.ACTIVE_LOW_BEGINTRANSFER       (1),
		.CHIPSELECT_THROUGH_READLATENCY (1)
	) ssram0 (
		.clk_clk                 (pcie_clk_clk),                               //   clk.clk
		.reset_reset             (rst_controller_001_reset_out_reset),         // reset.reset
		.uas_address             (mm_interconnect_0_ssram0_uas_address),       //   uas.address
		.uas_burstcount          (mm_interconnect_0_ssram0_uas_burstcount),    //      .burstcount
		.uas_read                (mm_interconnect_0_ssram0_uas_read),          //      .read
		.uas_write               (mm_interconnect_0_ssram0_uas_write),         //      .write
		.uas_waitrequest         (mm_interconnect_0_ssram0_uas_waitrequest),   //      .waitrequest
		.uas_readdatavalid       (mm_interconnect_0_ssram0_uas_readdatavalid), //      .readdatavalid
		.uas_byteenable          (mm_interconnect_0_ssram0_uas_byteenable),    //      .byteenable
		.uas_readdata            (mm_interconnect_0_ssram0_uas_readdata),      //      .readdata
		.uas_writedata           (mm_interconnect_0_ssram0_uas_writedata),     //      .writedata
		.uas_lock                (mm_interconnect_0_ssram0_uas_lock),          //      .lock
		.uas_debugaccess         (mm_interconnect_0_ssram0_uas_debugaccess),   //      .debugaccess
		.tcm_write_n_out         (ssram0_tcm_write_n_out),                     //   tcm.write_n_out
		.tcm_begintransfer_n_out (ssram0_tcm_begintransfer_n_out),             //      .begintransfer_n_out
		.tcm_chipselect_n_out    (ssram0_tcm_chipselect_n_out),                //      .chipselect_n_out
		.tcm_outputenable_n_out  (ssram0_tcm_outputenable_n_out),              //      .outputenable_n_out
		.tcm_request             (ssram0_tcm_request),                         //      .request
		.tcm_grant               (ssram0_tcm_grant),                           //      .grant
		.tcm_address_out         (ssram0_tcm_address_out),                     //      .address_out
		.tcm_byteenable_n_out    (ssram0_tcm_byteenable_n_out),                //      .byteenable_n_out
		.tcm_data_out            (ssram0_tcm_data_out),                        //      .data_out
		.tcm_data_outen          (ssram0_tcm_data_outen),                      //      .data_outen
		.tcm_data_in             (ssram0_tcm_data_in)                          //      .data_in
	);

	de2i_150_qsys_ssram0 #(
		.TCM_ADDRESS_W                  (22),
		.TCM_DATA_W                     (32),
		.TCM_BYTEENABLE_W               (4),
		.TCM_READ_WAIT                  (0),
		.TCM_WRITE_WAIT                 (0),
		.TCM_SETUP_WAIT                 (0),
		.TCM_DATA_HOLD                  (0),
		.TCM_TURNAROUND_TIME            (2),
		.TCM_TIMING_UNITS               (1),
		.TCM_READLATENCY                (4),
		.TCM_SYMBOLS_PER_WORD           (4),
		.USE_READDATA                   (1),
		.USE_WRITEDATA                  (1),
		.USE_READ                       (0),
		.USE_WRITE                      (1),
		.USE_BYTEENABLE                 (1),
		.USE_CHIPSELECT                 (1),
		.USE_LOCK                       (0),
		.USE_ADDRESS                    (1),
		.USE_WAITREQUEST                (0),
		.USE_WRITEBYTEENABLE            (0),
		.USE_OUTPUTENABLE               (1),
		.USE_RESETREQUEST               (0),
		.USE_IRQ                        (0),
		.USE_RESET_OUTPUT               (0),
		.ACTIVE_LOW_READ                (0),
		.ACTIVE_LOW_LOCK                (0),
		.ACTIVE_LOW_WRITE               (1),
		.ACTIVE_LOW_CHIPSELECT          (1),
		.ACTIVE_LOW_BYTEENABLE          (1),
		.ACTIVE_LOW_OUTPUTENABLE        (1),
		.ACTIVE_LOW_WRITEBYTEENABLE     (0),
		.ACTIVE_LOW_WAITREQUEST         (0),
		.ACTIVE_LOW_BEGINTRANSFER       (1),
		.CHIPSELECT_THROUGH_READLATENCY (1)
	) ssram1 (
		.clk_clk                 (pcie_clk_clk),                               //   clk.clk
		.reset_reset             (rst_controller_001_reset_out_reset),         // reset.reset
		.uas_address             (mm_interconnect_0_ssram1_uas_address),       //   uas.address
		.uas_burstcount          (mm_interconnect_0_ssram1_uas_burstcount),    //      .burstcount
		.uas_read                (mm_interconnect_0_ssram1_uas_read),          //      .read
		.uas_write               (mm_interconnect_0_ssram1_uas_write),         //      .write
		.uas_waitrequest         (mm_interconnect_0_ssram1_uas_waitrequest),   //      .waitrequest
		.uas_readdatavalid       (mm_interconnect_0_ssram1_uas_readdatavalid), //      .readdatavalid
		.uas_byteenable          (mm_interconnect_0_ssram1_uas_byteenable),    //      .byteenable
		.uas_readdata            (mm_interconnect_0_ssram1_uas_readdata),      //      .readdata
		.uas_writedata           (mm_interconnect_0_ssram1_uas_writedata),     //      .writedata
		.uas_lock                (mm_interconnect_0_ssram1_uas_lock),          //      .lock
		.uas_debugaccess         (mm_interconnect_0_ssram1_uas_debugaccess),   //      .debugaccess
		.tcm_write_n_out         (ssram1_tcm_write_n_out),                     //   tcm.write_n_out
		.tcm_begintransfer_n_out (ssram1_tcm_begintransfer_n_out),             //      .begintransfer_n_out
		.tcm_chipselect_n_out    (ssram1_tcm_chipselect_n_out),                //      .chipselect_n_out
		.tcm_outputenable_n_out  (ssram1_tcm_outputenable_n_out),              //      .outputenable_n_out
		.tcm_request             (ssram1_tcm_request),                         //      .request
		.tcm_grant               (ssram1_tcm_grant),                           //      .grant
		.tcm_address_out         (ssram1_tcm_address_out),                     //      .address_out
		.tcm_byteenable_n_out    (ssram1_tcm_byteenable_n_out),                //      .byteenable_n_out
		.tcm_data_out            (ssram1_tcm_data_out),                        //      .data_out
		.tcm_data_outen          (ssram1_tcm_data_outen),                      //      .data_outen
		.tcm_data_in             (ssram1_tcm_data_in)                          //      .data_in
	);

	de2i_150_qsys_tristate_conduit_bridge_0 tristate_conduit_bridge_0 (
		.clk               (pcie_clk_clk),                                       //   clk.clk
		.reset             (rst_controller_001_reset_out_reset),                 // reset.reset
		.request           (tristate_conduit_pin_sharer_0_tcm_request),          //   tcs.request
		.grant             (tristate_conduit_pin_sharer_0_tcm_grant),            //      .grant
		.tcs_ssram1_cs_n   (tristate_conduit_pin_sharer_0_tcm_ssram1_cs_n_out),  //      .ssram1_cs_n_out
		.tcs_ssram_adsc_n  (tristate_conduit_pin_sharer_0_tcm_ssram_adsc_n_out), //      .ssram_adsc_n_out
		.tcs_ssram_we_n    (tristate_conduit_pin_sharer_0_tcm_ssram_we_n_out),   //      .ssram_we_n_out
		.tcs_ssram_oe_n    (tristate_conduit_pin_sharer_0_tcm_ssram_oe_n_out),   //      .ssram_oe_n_out
		.tcs_fs_data       (tristate_conduit_pin_sharer_0_tcm_fs_data_out),      //      .fs_data_out
		.tcs_fs_data_outen (tristate_conduit_pin_sharer_0_tcm_fs_data_outen),    //      .fs_data_outen
		.tcs_fs_data_in    (tristate_conduit_pin_sharer_0_tcm_fs_data_in),       //      .fs_data_in
		.tcs_ssram_be_n    (tristate_conduit_pin_sharer_0_tcm_ssram_be_n_out),   //      .ssram_be_n_out
		.tcs_ssram0_cs_n   (tristate_conduit_pin_sharer_0_tcm_ssram0_cs_n_out),  //      .ssram0_cs_n_out
		.tcs_fs_addr       (tristate_conduit_pin_sharer_0_tcm_fs_addr_out),      //      .fs_addr_out
		.ssram1_cs_n       (flash_ssram_tri_state_bridge_out_ssram1_cs_n),       //   out.ssram1_cs_n
		.ssram_adsc_n      (flash_ssram_tri_state_bridge_out_ssram_adsc_n),      //      .ssram_adsc_n
		.ssram_we_n        (flash_ssram_tri_state_bridge_out_ssram_we_n),        //      .ssram_we_n
		.ssram_oe_n        (flash_ssram_tri_state_bridge_out_ssram_oe_n),        //      .ssram_oe_n
		.fs_data           (flash_ssram_tri_state_bridge_out_fs_data),           //      .fs_data
		.ssram_be_n        (flash_ssram_tri_state_bridge_out_ssram_be_n),        //      .ssram_be_n
		.ssram0_cs_n       (flash_ssram_tri_state_bridge_out_ssram0_cs_n),       //      .ssram0_cs_n
		.fs_addr           (flash_ssram_tri_state_bridge_out_fs_addr)            //      .fs_addr
	);

	de2i_150_qsys_tristate_conduit_pin_sharer_0 tristate_conduit_pin_sharer_0 (
		.clk_clk                  (pcie_clk_clk),                                       //   clk.clk
		.reset_reset              (rst_controller_001_reset_out_reset),                 // reset.reset
		.request                  (tristate_conduit_pin_sharer_0_tcm_request),          //   tcm.request
		.grant                    (tristate_conduit_pin_sharer_0_tcm_grant),            //      .grant
		.ssram1_cs_n              (tristate_conduit_pin_sharer_0_tcm_ssram1_cs_n_out),  //      .ssram1_cs_n_out
		.fs_addr                  (tristate_conduit_pin_sharer_0_tcm_fs_addr_out),      //      .fs_addr_out
		.ssram_be_n               (tristate_conduit_pin_sharer_0_tcm_ssram_be_n_out),   //      .ssram_be_n_out
		.ssram_oe_n               (tristate_conduit_pin_sharer_0_tcm_ssram_oe_n_out),   //      .ssram_oe_n_out
		.ssram_adsc_n             (tristate_conduit_pin_sharer_0_tcm_ssram_adsc_n_out), //      .ssram_adsc_n_out
		.ssram_we_n               (tristate_conduit_pin_sharer_0_tcm_ssram_we_n_out),   //      .ssram_we_n_out
		.fs_data                  (tristate_conduit_pin_sharer_0_tcm_fs_data_out),      //      .fs_data_out
		.fs_data_in               (tristate_conduit_pin_sharer_0_tcm_fs_data_in),       //      .fs_data_in
		.fs_data_outen            (tristate_conduit_pin_sharer_0_tcm_fs_data_outen),    //      .fs_data_outen
		.ssram0_cs_n              (tristate_conduit_pin_sharer_0_tcm_ssram0_cs_n_out),  //      .ssram0_cs_n_out
		.tcs0_request             (ssram0_tcm_request),                                 //  tcs0.request
		.tcs0_grant               (ssram0_tcm_grant),                                   //      .grant
		.tcs0_address_out         (ssram0_tcm_address_out),                             //      .address_out
		.tcs0_byteenable_n_out    (ssram0_tcm_byteenable_n_out),                        //      .byteenable_n_out
		.tcs0_outputenable_n_out  (ssram0_tcm_outputenable_n_out),                      //      .outputenable_n_out
		.tcs0_begintransfer_n_out (ssram0_tcm_begintransfer_n_out),                     //      .begintransfer_n_out
		.tcs0_write_n_out         (ssram0_tcm_write_n_out),                             //      .write_n_out
		.tcs0_data_out            (ssram0_tcm_data_out),                                //      .data_out
		.tcs0_data_in             (ssram0_tcm_data_in),                                 //      .data_in
		.tcs0_data_outen          (ssram0_tcm_data_outen),                              //      .data_outen
		.tcs0_chipselect_n_out    (ssram0_tcm_chipselect_n_out),                        //      .chipselect_n_out
		.tcs1_request             (ssram1_tcm_request),                                 //  tcs1.request
		.tcs1_grant               (ssram1_tcm_grant),                                   //      .grant
		.tcs1_address_out         (ssram1_tcm_address_out),                             //      .address_out
		.tcs1_byteenable_n_out    (ssram1_tcm_byteenable_n_out),                        //      .byteenable_n_out
		.tcs1_outputenable_n_out  (ssram1_tcm_outputenable_n_out),                      //      .outputenable_n_out
		.tcs1_begintransfer_n_out (ssram1_tcm_begintransfer_n_out),                     //      .begintransfer_n_out
		.tcs1_write_n_out         (ssram1_tcm_write_n_out),                             //      .write_n_out
		.tcs1_data_out            (ssram1_tcm_data_out),                                //      .data_out
		.tcs1_data_in             (ssram1_tcm_data_in),                                 //      .data_in
		.tcs1_data_outen          (ssram1_tcm_data_outen),                              //      .data_outen
		.tcs1_chipselect_n_out    (ssram1_tcm_chipselect_n_out)                         //      .chipselect_n_out
	);

	de2i_150_qsys_height width (
		.clk      (pcie_clk_clk),                        //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset), //               reset.reset_n
		.address  (mm_interconnect_0_width_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_width_s1_readdata), //                    .readdata
		.in_port  (width_external_connection_export)     // external_connection.export
	);

	de2i_150_qsys_mm_interconnect_0 mm_interconnect_0 (
		.altpll_0_c1_clk                                             (altpll_0_c1_clk),                               //                                           altpll_0_c1.clk
		.pcie_ip_pcie_core_clk_clk                                   (pcie_clk_clk),                                  //                                 pcie_ip_pcie_core_clk.clk
		.mem_master_clock_reset_reset_reset_bridge_in_reset_reset    (rst_controller_001_reset_out_reset),            //    mem_master_clock_reset_reset_reset_bridge_in_reset.reset
		.pcie_ip_bar1_0_translator_reset_reset_bridge_in_reset_reset (rst_controller_003_reset_out_reset),            // pcie_ip_bar1_0_translator_reset_reset_bridge_in_reset.reset
		.sram0_reset_reset_bridge_in_reset_reset                     (rst_controller_002_reset_out_reset),            //                     sram0_reset_reset_bridge_in_reset.reset
		.mem_master_avalon_master_address                            (mem_master_avalon_master_address),              //                              mem_master_avalon_master.address
		.mem_master_avalon_master_waitrequest                        (mem_master_avalon_master_waitrequest),          //                                                      .waitrequest
		.mem_master_avalon_master_burstcount                         (mem_master_avalon_master_burstcount),           //                                                      .burstcount
		.mem_master_avalon_master_byteenable                         (mem_master_avalon_master_byteenable),           //                                                      .byteenable
		.mem_master_avalon_master_read                               (mem_master_avalon_master_read),                 //                                                      .read
		.mem_master_avalon_master_readdata                           (mem_master_avalon_master_readdata),             //                                                      .readdata
		.mem_master_avalon_master_readdatavalid                      (mem_master_avalon_master_readdatavalid),        //                                                      .readdatavalid
		.pcie_ip_bar1_0_address                                      (pcie_ip_bar1_0_address),                        //                                        pcie_ip_bar1_0.address
		.pcie_ip_bar1_0_waitrequest                                  (pcie_ip_bar1_0_waitrequest),                    //                                                      .waitrequest
		.pcie_ip_bar1_0_burstcount                                   (pcie_ip_bar1_0_burstcount),                     //                                                      .burstcount
		.pcie_ip_bar1_0_byteenable                                   (pcie_ip_bar1_0_byteenable),                     //                                                      .byteenable
		.pcie_ip_bar1_0_read                                         (pcie_ip_bar1_0_read),                           //                                                      .read
		.pcie_ip_bar1_0_readdata                                     (pcie_ip_bar1_0_readdata),                       //                                                      .readdata
		.pcie_ip_bar1_0_readdatavalid                                (pcie_ip_bar1_0_readdatavalid),                  //                                                      .readdatavalid
		.pcie_ip_bar1_0_write                                        (pcie_ip_bar1_0_write),                          //                                                      .write
		.pcie_ip_bar1_0_writedata                                    (pcie_ip_bar1_0_writedata),                      //                                                      .writedata
		.sgdma_descriptor_read_address                               (sgdma_descriptor_read_address),                 //                                 sgdma_descriptor_read.address
		.sgdma_descriptor_read_waitrequest                           (sgdma_descriptor_read_waitrequest),             //                                                      .waitrequest
		.sgdma_descriptor_read_read                                  (sgdma_descriptor_read_read),                    //                                                      .read
		.sgdma_descriptor_read_readdata                              (sgdma_descriptor_read_readdata),                //                                                      .readdata
		.sgdma_descriptor_read_readdatavalid                         (sgdma_descriptor_read_readdatavalid),           //                                                      .readdatavalid
		.sgdma_descriptor_write_address                              (sgdma_descriptor_write_address),                //                                sgdma_descriptor_write.address
		.sgdma_descriptor_write_waitrequest                          (sgdma_descriptor_write_waitrequest),            //                                                      .waitrequest
		.sgdma_descriptor_write_write                                (sgdma_descriptor_write_write),                  //                                                      .write
		.sgdma_descriptor_write_writedata                            (sgdma_descriptor_write_writedata),              //                                                      .writedata
		.sgdma_m_read_address                                        (sgdma_m_read_address),                          //                                          sgdma_m_read.address
		.sgdma_m_read_waitrequest                                    (sgdma_m_read_waitrequest),                      //                                                      .waitrequest
		.sgdma_m_read_read                                           (sgdma_m_read_read),                             //                                                      .read
		.sgdma_m_read_readdata                                       (sgdma_m_read_readdata),                         //                                                      .readdata
		.sgdma_m_read_readdatavalid                                  (sgdma_m_read_readdatavalid),                    //                                                      .readdatavalid
		.sgdma_m_write_address                                       (sgdma_m_write_address),                         //                                         sgdma_m_write.address
		.sgdma_m_write_waitrequest                                   (sgdma_m_write_waitrequest),                     //                                                      .waitrequest
		.sgdma_m_write_byteenable                                    (sgdma_m_write_byteenable),                      //                                                      .byteenable
		.sgdma_m_write_write                                         (sgdma_m_write_write),                           //                                                      .write
		.sgdma_m_write_writedata                                     (sgdma_m_write_writedata),                       //                                                      .writedata
		.button_s1_address                                           (mm_interconnect_0_button_s1_address),           //                                             button_s1.address
		.button_s1_write                                             (mm_interconnect_0_button_s1_write),             //                                                      .write
		.button_s1_readdata                                          (mm_interconnect_0_button_s1_readdata),          //                                                      .readdata
		.button_s1_writedata                                         (mm_interconnect_0_button_s1_writedata),         //                                                      .writedata
		.button_s1_chipselect                                        (mm_interconnect_0_button_s1_chipselect),        //                                                      .chipselect
		.chip_sel_s1_address                                         (mm_interconnect_0_chip_sel_s1_address),         //                                           chip_sel_s1.address
		.chip_sel_s1_write                                           (mm_interconnect_0_chip_sel_s1_write),           //                                                      .write
		.chip_sel_s1_readdata                                        (mm_interconnect_0_chip_sel_s1_readdata),        //                                                      .readdata
		.chip_sel_s1_writedata                                       (mm_interconnect_0_chip_sel_s1_writedata),       //                                                      .writedata
		.chip_sel_s1_chipselect                                      (mm_interconnect_0_chip_sel_s1_chipselect),      //                                                      .chipselect
		.height_s1_address                                           (mm_interconnect_0_height_s1_address),           //                                             height_s1.address
		.height_s1_readdata                                          (mm_interconnect_0_height_s1_readdata),          //                                                      .readdata
		.led_s1_address                                              (mm_interconnect_0_led_s1_address),              //                                                led_s1.address
		.led_s1_write                                                (mm_interconnect_0_led_s1_write),                //                                                      .write
		.led_s1_readdata                                             (mm_interconnect_0_led_s1_readdata),             //                                                      .readdata
		.led_s1_writedata                                            (mm_interconnect_0_led_s1_writedata),            //                                                      .writedata
		.led_s1_chipselect                                           (mm_interconnect_0_led_s1_chipselect),           //                                                      .chipselect
		.onchip_memory_s1_address                                    (mm_interconnect_0_onchip_memory_s1_address),    //                                      onchip_memory_s1.address
		.onchip_memory_s1_write                                      (mm_interconnect_0_onchip_memory_s1_write),      //                                                      .write
		.onchip_memory_s1_readdata                                   (mm_interconnect_0_onchip_memory_s1_readdata),   //                                                      .readdata
		.onchip_memory_s1_writedata                                  (mm_interconnect_0_onchip_memory_s1_writedata),  //                                                      .writedata
		.onchip_memory_s1_byteenable                                 (mm_interconnect_0_onchip_memory_s1_byteenable), //                                                      .byteenable
		.onchip_memory_s1_chipselect                                 (mm_interconnect_0_onchip_memory_s1_chipselect), //                                                      .chipselect
		.onchip_memory_s1_clken                                      (mm_interconnect_0_onchip_memory_s1_clken),      //                                                      .clken
		.pcie_ip_txs_address                                         (mm_interconnect_0_pcie_ip_txs_address),         //                                           pcie_ip_txs.address
		.pcie_ip_txs_write                                           (mm_interconnect_0_pcie_ip_txs_write),           //                                                      .write
		.pcie_ip_txs_read                                            (mm_interconnect_0_pcie_ip_txs_read),            //                                                      .read
		.pcie_ip_txs_readdata                                        (mm_interconnect_0_pcie_ip_txs_readdata),        //                                                      .readdata
		.pcie_ip_txs_writedata                                       (mm_interconnect_0_pcie_ip_txs_writedata),       //                                                      .writedata
		.pcie_ip_txs_burstcount                                      (mm_interconnect_0_pcie_ip_txs_burstcount),      //                                                      .burstcount
		.pcie_ip_txs_byteenable                                      (mm_interconnect_0_pcie_ip_txs_byteenable),      //                                                      .byteenable
		.pcie_ip_txs_readdatavalid                                   (mm_interconnect_0_pcie_ip_txs_readdatavalid),   //                                                      .readdatavalid
		.pcie_ip_txs_waitrequest                                     (mm_interconnect_0_pcie_ip_txs_waitrequest),     //                                                      .waitrequest
		.pcie_ip_txs_chipselect                                      (mm_interconnect_0_pcie_ip_txs_chipselect),      //                                                      .chipselect
		.pio_size_s1_address                                         (mm_interconnect_0_pio_size_s1_address),         //                                           pio_size_s1.address
		.pio_size_s1_write                                           (mm_interconnect_0_pio_size_s1_write),           //                                                      .write
		.pio_size_s1_readdata                                        (mm_interconnect_0_pio_size_s1_readdata),        //                                                      .readdata
		.pio_size_s1_writedata                                       (mm_interconnect_0_pio_size_s1_writedata),       //                                                      .writedata
		.pio_size_s1_chipselect                                      (mm_interconnect_0_pio_size_s1_chipselect),      //                                                      .chipselect
		.sram0_s1_address                                            (mm_interconnect_0_sram0_s1_address),            //                                              sram0_s1.address
		.sram0_s1_write                                              (mm_interconnect_0_sram0_s1_write),              //                                                      .write
		.sram0_s1_read                                               (mm_interconnect_0_sram0_s1_read),               //                                                      .read
		.sram0_s1_readdata                                           (mm_interconnect_0_sram0_s1_readdata),           //                                                      .readdata
		.sram0_s1_writedata                                          (mm_interconnect_0_sram0_s1_writedata),          //                                                      .writedata
		.sram0_s1_byteenable                                         (mm_interconnect_0_sram0_s1_byteenable),         //                                                      .byteenable
		.sram0_s1_readdatavalid                                      (mm_interconnect_0_sram0_s1_readdatavalid),      //                                                      .readdatavalid
		.sram0_s1_waitrequest                                        (mm_interconnect_0_sram0_s1_waitrequest),        //                                                      .waitrequest
		.sram0_s1_chipselect                                         (mm_interconnect_0_sram0_s1_chipselect),         //                                                      .chipselect
		.ssram0_uas_address                                          (mm_interconnect_0_ssram0_uas_address),          //                                            ssram0_uas.address
		.ssram0_uas_write                                            (mm_interconnect_0_ssram0_uas_write),            //                                                      .write
		.ssram0_uas_read                                             (mm_interconnect_0_ssram0_uas_read),             //                                                      .read
		.ssram0_uas_readdata                                         (mm_interconnect_0_ssram0_uas_readdata),         //                                                      .readdata
		.ssram0_uas_writedata                                        (mm_interconnect_0_ssram0_uas_writedata),        //                                                      .writedata
		.ssram0_uas_burstcount                                       (mm_interconnect_0_ssram0_uas_burstcount),       //                                                      .burstcount
		.ssram0_uas_byteenable                                       (mm_interconnect_0_ssram0_uas_byteenable),       //                                                      .byteenable
		.ssram0_uas_readdatavalid                                    (mm_interconnect_0_ssram0_uas_readdatavalid),    //                                                      .readdatavalid
		.ssram0_uas_waitrequest                                      (mm_interconnect_0_ssram0_uas_waitrequest),      //                                                      .waitrequest
		.ssram0_uas_lock                                             (mm_interconnect_0_ssram0_uas_lock),             //                                                      .lock
		.ssram0_uas_debugaccess                                      (mm_interconnect_0_ssram0_uas_debugaccess),      //                                                      .debugaccess
		.ssram1_uas_address                                          (mm_interconnect_0_ssram1_uas_address),          //                                            ssram1_uas.address
		.ssram1_uas_write                                            (mm_interconnect_0_ssram1_uas_write),            //                                                      .write
		.ssram1_uas_read                                             (mm_interconnect_0_ssram1_uas_read),             //                                                      .read
		.ssram1_uas_readdata                                         (mm_interconnect_0_ssram1_uas_readdata),         //                                                      .readdata
		.ssram1_uas_writedata                                        (mm_interconnect_0_ssram1_uas_writedata),        //                                                      .writedata
		.ssram1_uas_burstcount                                       (mm_interconnect_0_ssram1_uas_burstcount),       //                                                      .burstcount
		.ssram1_uas_byteenable                                       (mm_interconnect_0_ssram1_uas_byteenable),       //                                                      .byteenable
		.ssram1_uas_readdatavalid                                    (mm_interconnect_0_ssram1_uas_readdatavalid),    //                                                      .readdatavalid
		.ssram1_uas_waitrequest                                      (mm_interconnect_0_ssram1_uas_waitrequest),      //                                                      .waitrequest
		.ssram1_uas_lock                                             (mm_interconnect_0_ssram1_uas_lock),             //                                                      .lock
		.ssram1_uas_debugaccess                                      (mm_interconnect_0_ssram1_uas_debugaccess),      //                                                      .debugaccess
		.width_s1_address                                            (mm_interconnect_0_width_s1_address),            //                                              width_s1.address
		.width_s1_readdata                                           (mm_interconnect_0_width_s1_readdata)            //                                                      .readdata
	);

	de2i_150_qsys_mm_interconnect_1 mm_interconnect_1 (
		.pcie_ip_pcie_core_clk_clk                                 (pcie_clk_clk),                              //                               pcie_ip_pcie_core_clk.clk
		.pcie_ip_bar2_translator_reset_reset_bridge_in_reset_reset (rst_controller_003_reset_out_reset),        // pcie_ip_bar2_translator_reset_reset_bridge_in_reset.reset
		.sgdma_reset_reset_bridge_in_reset_reset                   (rst_controller_001_reset_out_reset),        //                   sgdma_reset_reset_bridge_in_reset.reset
		.pcie_ip_bar2_address                                      (pcie_ip_bar2_address),                      //                                        pcie_ip_bar2.address
		.pcie_ip_bar2_waitrequest                                  (pcie_ip_bar2_waitrequest),                  //                                                    .waitrequest
		.pcie_ip_bar2_burstcount                                   (pcie_ip_bar2_burstcount),                   //                                                    .burstcount
		.pcie_ip_bar2_byteenable                                   (pcie_ip_bar2_byteenable),                   //                                                    .byteenable
		.pcie_ip_bar2_read                                         (pcie_ip_bar2_read),                         //                                                    .read
		.pcie_ip_bar2_readdata                                     (pcie_ip_bar2_readdata),                     //                                                    .readdata
		.pcie_ip_bar2_readdatavalid                                (pcie_ip_bar2_readdatavalid),                //                                                    .readdatavalid
		.pcie_ip_bar2_write                                        (pcie_ip_bar2_write),                        //                                                    .write
		.pcie_ip_bar2_writedata                                    (pcie_ip_bar2_writedata),                    //                                                    .writedata
		.pcie_ip_cra_address                                       (mm_interconnect_1_pcie_ip_cra_address),     //                                         pcie_ip_cra.address
		.pcie_ip_cra_write                                         (mm_interconnect_1_pcie_ip_cra_write),       //                                                    .write
		.pcie_ip_cra_read                                          (mm_interconnect_1_pcie_ip_cra_read),        //                                                    .read
		.pcie_ip_cra_readdata                                      (mm_interconnect_1_pcie_ip_cra_readdata),    //                                                    .readdata
		.pcie_ip_cra_writedata                                     (mm_interconnect_1_pcie_ip_cra_writedata),   //                                                    .writedata
		.pcie_ip_cra_byteenable                                    (mm_interconnect_1_pcie_ip_cra_byteenable),  //                                                    .byteenable
		.pcie_ip_cra_waitrequest                                   (mm_interconnect_1_pcie_ip_cra_waitrequest), //                                                    .waitrequest
		.pcie_ip_cra_chipselect                                    (mm_interconnect_1_pcie_ip_cra_chipselect),  //                                                    .chipselect
		.sgdma_csr_address                                         (mm_interconnect_1_sgdma_csr_address),       //                                           sgdma_csr.address
		.sgdma_csr_write                                           (mm_interconnect_1_sgdma_csr_write),         //                                                    .write
		.sgdma_csr_read                                            (mm_interconnect_1_sgdma_csr_read),          //                                                    .read
		.sgdma_csr_readdata                                        (mm_interconnect_1_sgdma_csr_readdata),      //                                                    .readdata
		.sgdma_csr_writedata                                       (mm_interconnect_1_sgdma_csr_writedata),     //                                                    .writedata
		.sgdma_csr_chipselect                                      (mm_interconnect_1_sgdma_csr_chipselect)     //                                                    .chipselect
	);

	de2i_150_qsys_irq_mapper irq_mapper (
		.clk           (pcie_clk_clk),                       //       clk.clk
		.reset         (rst_controller_003_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.sender_irq    (pcie_ip_rxm_irq_irq)                 //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.reset_in1      (~pcie_ip_pcie_core_reset_reset), // reset_in1.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (~pcie_ip_pcie_core_reset_reset),         // reset_in1.reset
		.clk            (pcie_clk_clk),                           //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (~pcie_ip_pcie_core_reset_reset),     // reset_in1.reset
		.clk            (altpll_0_c1_clk),                    //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_003 (
		.reset_in0      (~pcie_ip_pcie_core_reset_reset),     // reset_in0.reset
		.clk            (pcie_clk_clk),                       //       clk.clk
		.reset_out      (rst_controller_003_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	assign pcie_rst_n_reset_n = ~rst_controller_001_reset_out_reset;

endmodule
